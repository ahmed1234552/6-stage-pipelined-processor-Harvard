LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
entity controller is
    port (
      opcode : in std_logic_vector(4 downto 0);
      wb : out std_logic ;
      mem_rd : out std_logic;
      mem_wr : out std_logic;
      stck_wr : out std_logic;
      stck_rd : out std_logic;
      pc_to_stck : out std_logic;
      port_wr : out std_logic;
      port_rd : out std_logic;
      ldm : out std_logic;
      alu_op : out std_logic; -- it could be 2 bits
      rtrn_pc_signal : out std_logic;
      rti : out std_logic;
      alu_src : out std_logic;
      branch : out std_logic
    );
end entity;

architecture behavioral of controller is
  begin
    process (opcode)
    begin
      case opcode is
        when "00000" => -- NOP
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0';
          branch <= '0';
        when "00001" => -- Clrc
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0';
          branch <= '0';
        when "00010" => -- setc
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0';
          branch <= '0';
        when "00011" => -- Dec
          wb <= '1';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "00100" => -- Inc
          wb <= '1';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "00101" => -- Out
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '1';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "00110" => -- In
          wb <= '1';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '1';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0'; ----------------------------------------------------------------
        when "01000" => -- mov 
          wb <= '1';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "01001" => -- Not 
          wb <= '1';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0'; 
        when "01010" => -- Add 
          wb <= '1';
          mem_rd <= '0'; -- 0 for read, 1 for write
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '1'; 
          branch <= '0';
        when "01011" => -- Sub 
          wb <= '1';
          mem_rd <= '0'; -- 0 for read, 1 for write
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '1'; 
          branch <= '0';
        when "01100" => -- AND 
          wb <= '1';
          mem_rd <= '0'; -- 0 for read, 1 for write
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '1'; 
          branch <= '0';
        when "01101" => -- OR 
          wb <= '1';
          mem_rd <= '0'; -- 0 for read, 1 for write
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '1'; 
          branch <= '0';
        when "01110" => -- IADD 
          wb <= '1';
          mem_rd <= '0'; -- 0 for read, 1 for write
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '1';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; 
          branch <= '0'; ----------------------------------------------------------------
        when "10000" => -- PUSH 
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '1';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "10001" => -- POP 
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '1';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "10010" => -- LDM 
          wb <= '1';
          mem_rd <= '1';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '1';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "10011" => -- LDD 1	1	0	0	0	0	0	0	0	0	0	0	X	0
          wb <= '1';
          mem_rd <= '1';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "10100" => -- STD 0	0	1	0	0	0	0	0	0	0	0	0	X	0
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '1';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0'; ----------------------------------------------------------------
        when "11000" => -- JZ 
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '1';
        when "11001" => -- JN -- JNZ  
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '1';
        when "11010" => -- JC 
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '1';
        when "11011" => -- JMP 
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "11100" => -- CALL 0	0	0	1	0	1	0	0	0	0	0	0	X	0
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '1';
          stck_rd <= '0';
          pc_to_stck <= '1';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "11101" => -- RET 0	0	0	0	1	0	0	0	0	0	1	0	X	0
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '1';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '1';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when "11110" => -- RTI 0	0	0	0	1	0	0	0	0	0	1	1	X	0
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '1';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '1';
          rti <= '1';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
        when others =>
          wb <= '0';
          mem_rd <= '0';
          mem_wr <= '0';
          stck_wr <= '0';
          stck_rd <= '0';
          pc_to_stck <= '0';
          port_wr <= '0';
          port_rd <= '0';
          ldm <= '0';
          alu_op <= '0';
          rtrn_pc_signal <= '0';
          rti <= '0';
          alu_src <= '0'; -- 0 for A, 1 for B
          branch <= '0';
      end case;
    end process;
end architecture behavioral;


        

          
          
          
          
